module fsm (
    input        clk,
    input        rst,
    output [4:0] leds,     // flag LEDs
    output [3:0] bcd_out,  // BCD to show
    output       buzzer    // buzzer signal
);

endmodule  //fsm

//-----------------------------------------------------------------------------
//
// Title       : calc
// Design      : calc
// Author      : aheir
// Company     : aheir
//
//-----------------------------------------------------------------------------
//
// File        : F:\documents\alheir\e3-2022-tp2\active\e3tp2\src\calc.v
// Generated   : Sun Oct 30 22:02:15 2022
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {calc}}
module calc ();

//}} End of automatically maintained section

// -- Enter your statements here -- //

endmodule

module display (
    input clk,
    input rst,
    input [3:0] a  // BCD to show
);

endmodule  //display
